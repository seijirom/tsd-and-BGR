* Created by KLayout

* cell bgr8
* pin R1
* pin R3
* pin R2
* pin SUBSTRATE
.SUBCKT bgr8 3 14 23 35
* net 3 R1
* net 14 R3
* net 23 R2
* net 35 SUBSTRATE
* device instance $3 r0 *1 -45,-108.5 RES
R$3 4 1 4000 RES
* device instance $18 m0 *1 171,-96.5 RES
R$18 23 3 4000 RES
* device instance $53 r0 *1 101,-184.5 RES
R$53 6 3 24000 RES
* device instance $58 m90 *1 -44.5,-199.5 RES
R$58 35 4 26000 RES
* device instance $73 r0 *1 90,-96.5 RES
R$73 13 14 2000 RES
* device instance $83 m90 *1 132,-96.5 RES
R$83 14 23 2000 RES
* device instance $101 r180 *1 -37.5,-20 HRES
R$101 24 26 1001000 HRES
* device instance $107 m90 *1 75.5,-59.5 D
D$107 35 19 D A=4P P=8U
* device instance $108 r90 *1 63.5,-56 D
D$108 35 20 D A=4P P=8U
* device instance $109 r0 *1 28,-73.5 NMOS
M$109 5 18 19 35 NMOS L=1U W=80U AS=160P AD=160P PS=176U PD=176U
* device instance $113 r0 *1 35,-110.5 NMOS
M$113 9 18 20 35 NMOS L=1U W=80U AS=160P AD=160P PS=176U PD=176U
* device instance $117 r0 *1 -13,-108.5 NMOS
M$117 13 18 18 35 NMOS L=1U W=160U AS=320P AD=320P PS=352U PD=352U
* device instance $125 r0 *1 91.5,-32.5 PMOS
M$125 34 19 18 24 PMOS L=1U W=20U AS=40P AD=40P PS=44U PD=44U
* device instance $126 r0 *1 63.5,-32.5 PMOS
M$126 32 19 18 24 PMOS L=1U W=20U AS=40P AD=40P PS=44U PD=44U
* device instance $127 r0 *1 49.5,-32.5 PMOS
M$127 31 19 18 24 PMOS L=1U W=20U AS=40P AD=40P PS=44U PD=44U
* device instance $128 r0 *1 77.5,-32.5 PMOS
M$128 33 19 18 24 PMOS L=1U W=20U AS=40P AD=40P PS=44U PD=44U
* device instance $129 r0 *1 35.5,-32 PMOS
M$129 30 19 19 24 PMOS L=1U W=20U AS=40P AD=40P PS=44U PD=44U
* device instance $130 r0 *1 88.5,2 PMOS
M$130 24 19 34 24 PMOS L=1U W=20U AS=40P AD=40P PS=44U PD=44U
* device instance $131 r0 *1 74.5,2 PMOS
M$131 24 19 33 24 PMOS L=1U W=20U AS=40P AD=40P PS=44U PD=44U
* device instance $132 r0 *1 32.5,2 PMOS
M$132 24 19 30 24 PMOS L=1U W=20U AS=40P AD=40P PS=44U PD=44U
* device instance $133 r0 *1 60.5,2 PMOS
M$133 24 19 32 24 PMOS L=1U W=20U AS=40P AD=40P PS=44U PD=44U
* device instance $134 r0 *1 46.5,2 PMOS
M$134 24 19 31 24 PMOS L=1U W=20U AS=40P AD=40P PS=44U PD=44U
* device instance $135 r0 *1 4.5,2 PMOS
M$135 24 19 28 24 PMOS L=1U W=20U AS=40P AD=40P PS=44U PD=44U
* device instance $136 r0 *1 7.5,-31.5 PMOS
M$136 28 19 20 24 PMOS L=1U W=20U AS=40P AD=40P PS=44U PD=44U
* device instance $137 r0 *1 21.5,-32 PMOS
M$137 29 20 19 24 PMOS L=1U W=20U AS=40P AD=40P PS=44U PD=44U
* device instance $138 r0 *1 -6.5,-32 PMOS
M$138 27 20 20 24 PMOS L=1U W=20U AS=40P AD=40P PS=44U PD=44U
* device instance $139 r0 *1 -9.5,2 PMOS
M$139 24 20 27 24 PMOS L=1U W=20U AS=40P AD=40P PS=44U PD=44U
* device instance $140 r0 *1 18.5,2 PMOS
M$140 24 20 29 24 PMOS L=1U W=20U AS=40P AD=40P PS=44U PD=44U
* device instance $141 r180 *1 -4.5,-211.5 PMOS
M$141 5 5 5 1 PMOS L=1U W=160U AS=320P AD=320P PS=352U PD=352U
* device instance $149 r180 *1 10,-179.5 PMOS
M$149 9 9 9 4 PMOS L=1U W=20U AS=40P AD=40P PS=44U PD=44U
* device instance $150 r180 *1 43,-173.5 PMOS
M$150 6 6 6 35 PMOS L=1U W=40U AS=80P AD=80P PS=88U PD=88U
.ENDS bgr8
