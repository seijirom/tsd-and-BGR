* Created by KLayout

* cell external
* pin SUBSTRATE
* pin $1.R35k
* pin $1.A
* pin $1.D
* pin $1.VOUT
* pin $1.R3
* pin $1.R2
* pin $1.R1
* pin $1.R25k
* pin $1.R50k
* pin $1.R65k
* pin $1.R75k
* pin $1.TSD
* pin $1.res1meg
* pin $1.VDD
* pin $1.ext1meg
* pin $1.B
.SUBCKT external 2 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19
* net 2 SUBSTRATE
* net 4 $1.R35k
* net 5 $1.A
* net 6 $1.D
* net 7 $1.VOUT
* net 8 $1.R3
* net 9 $1.R2
* net 10 $1.R1
* net 11 $1.R25k
* net 12 $1.R50k
* net 13 $1.R65k
* net 14 $1.R75k
* net 15 $1.TSD
* net 16 $1.res1meg
* net 17 $1.VDD
* net 18 $1.ext1meg
* net 19 $1.B
* cell instance $2 r0 *1 -1,-0.5
X$2 5 15 19 17 1 2 2 1 3 tsd_2021
* cell instance $3 r0 *1 -1,0
X$3 6 10 7 8 18 3 9 16 2 bgr8
* device instance $1 r0 *1 284.5,-33 HRES
R$1 5 14 75000 HRES
* device instance $2 r0 *1 147,-15.5 HRES
R$2 5 11 25000 HRES
* device instance $3 r0 *1 245,-34 HRES
R$3 5 13 65000 HRES
* device instance $4 r0 *1 178.5,-16 HRES
R$4 5 4 35000 HRES
* device instance $5 r0 *1 212.5,-31.5 HRES
R$5 5 12 50000 HRES
.ENDS external

* cell tsd_2021
* pin 
* pin 
* pin 
* pin 
* pin 
* pin SUBSTRATE
* pin 
* pin 
* pin 
.SUBCKT tsd_2021 1 2 4 7 8 9 10 11 12
* net 9 SUBSTRATE
* device instance $1 r0 *1 186,-218 NMOS
M$1 9 6 3 9 NMOS L=1U W=200U AS=220P AD=220P PS=242U PD=242U
* device instance $11 r0 *1 286,-218 NMOS
M$11 9 6 8 9 NMOS L=1U W=100U AS=120P AD=120P PS=132U PD=132U
* device instance $16 r0 *1 266,-202.5 HRES
R$16 10 1 20000 HRES
* device instance $17 r90 *1 297.5,-185 HRES
R$17 1 11 100000 HRES
* device instance $20 m90 *1 206.5,-185.5 NMOS
M$20 9 3 2 9 NMOS L=1U W=200U AS=220P AD=220P PS=242U PD=242U
* device instance $30 r0 *1 266.5,-112.5 PMOS
M$30 7 12 16 7 PMOS L=1U W=20U AS=40P AD=40P PS=44U PD=44U
* device instance $31 r0 *1 200.5,-112.5 PMOS
M$31 7 12 20 7 PMOS L=1U W=20U AS=40P AD=40P PS=44U PD=44U
* device instance $32 r0 *1 209.5,-112.5 PMOS
M$32 7 12 19 7 PMOS L=1U W=20U AS=40P AD=40P PS=44U PD=44U
* device instance $33 r0 *1 222.5,-112.5 PMOS
M$33 7 12 18 7 PMOS L=1U W=20U AS=40P AD=40P PS=44U PD=44U
* device instance $34 r0 *1 231.5,-112.5 PMOS
M$34 7 12 17 7 PMOS L=1U W=20U AS=40P AD=40P PS=44U PD=44U
* device instance $35 r0 *1 244.5,-112.5 PMOS
M$35 7 12 14 7 PMOS L=1U W=20U AS=40P AD=40P PS=44U PD=44U
* device instance $36 r0 *1 253.5,-112.5 PMOS
M$36 7 12 15 7 PMOS L=1U W=20U AS=40P AD=40P PS=44U PD=44U
* device instance $37 r0 *1 275.5,-112.5 PMOS
M$37 7 12 13 7 PMOS L=1U W=20U AS=40P AD=40P PS=44U PD=44U
* device instance $38 r0 *1 235,-214 NMOS
M$38 9 23 23 9 NMOS L=1U W=20U AS=40P AD=40P PS=44U PD=44U
* device instance $39 m90 *1 226.5,-214 NMOS
M$39 9 23 6 9 NMOS L=1U W=20U AS=40P AD=40P PS=44U PD=44U
* device instance $40 r180 *1 249,-214 PMOS
M$40 4 4 4 9 PMOS L=1U W=20U AS=40P AD=40P PS=44U PD=44U
* device instance $41 r180 *1 278.5,-143.5 PMOS
M$41 1 12 13 7 PMOS L=1U W=20U AS=40P AD=40P PS=44U PD=44U
* device instance $42 r180 *1 203.5,-144 PMOS
M$42 3 12 20 7 PMOS L=1U W=20U AS=40P AD=40P PS=44U PD=44U
* device instance $43 r180 *1 212.5,-144 PMOS
M$43 3 12 19 7 PMOS L=1U W=20U AS=40P AD=40P PS=44U PD=44U
* device instance $44 r180 *1 225.5,-143.5 PMOS
M$44 5 12 18 7 PMOS L=1U W=20U AS=40P AD=40P PS=44U PD=44U
* device instance $45 r180 *1 234.5,-143.5 PMOS
M$45 5 12 17 7 PMOS L=1U W=20U AS=40P AD=40P PS=44U PD=44U
* device instance $46 r180 *1 247.5,-143.5 PMOS
M$46 4 12 14 7 PMOS L=1U W=20U AS=40P AD=40P PS=44U PD=44U
* device instance $47 r180 *1 256.5,-143.5 PMOS
M$47 4 12 15 7 PMOS L=1U W=20U AS=40P AD=40P PS=44U PD=44U
* device instance $48 r180 *1 269.5,-143.5 PMOS
M$48 1 12 16 7 PMOS L=1U W=20U AS=40P AD=40P PS=44U PD=44U
* device instance $49 m90 *1 236,-185 PMOS
M$49 5 4 23 5 PMOS L=1U W=20U AS=40P AD=40P PS=44U PD=44U
* device instance $50 r0 *1 222.5,-185 PMOS
M$50 5 1 6 5 PMOS L=1U W=20U AS=40P AD=40P PS=44U PD=44U
.ENDS tsd_2021

* cell bgr8
* pin D
* pin R1
* pin Vout
* pin R3
* pin ext1meg
* pin VBG
* pin R2
* pin res1meg
* pin SUBSTRATE
.SUBCKT bgr8 3 4 16 17 18 19 23 24 35
* net 3 D
* net 4 R1
* net 16 Vout
* net 17 R3
* net 18 ext1meg
* net 19 VBG
* net 23 R2
* net 24 res1meg
* net 35 SUBSTRATE
* device instance $3 r0 *1 -45,-108.5 RES
R$3 5 1 4000 RES
* device instance $23 m0 *1 171,-96.5 RES
R$23 23 4 4000 RES
* device instance $53 r0 *1 101,-184.5 RES
R$53 3 4 24000 RES
* device instance $58 m90 *1 -24.5,-199.5 RES
R$58 35 5 26000 RES
* device instance $73 r0 *1 110,-96.5 RES
R$73 16 17 2000 RES
* device instance $83 m90 *1 132,-96.5 RES
R$83 17 23 2000 RES
* device instance $101 r0 *1 88.5,2 PMOS
M$101 25 19 34 25 PMOS L=1U W=20U AS=40P AD=40P PS=44U PD=44U
* device instance $102 r0 *1 74.5,2 PMOS
M$102 25 19 33 25 PMOS L=1U W=20U AS=40P AD=40P PS=44U PD=44U
* device instance $103 r0 *1 32.5,2 PMOS
M$103 25 19 30 25 PMOS L=1U W=20U AS=40P AD=40P PS=44U PD=44U
* device instance $104 r0 *1 60.5,2 PMOS
M$104 25 19 32 25 PMOS L=1U W=20U AS=40P AD=40P PS=44U PD=44U
* device instance $105 r0 *1 46.5,2 PMOS
M$105 25 19 31 25 PMOS L=1U W=20U AS=40P AD=40P PS=44U PD=44U
* device instance $106 r0 *1 4.5,2 PMOS
M$106 25 19 28 25 PMOS L=1U W=20U AS=40P AD=40P PS=44U PD=44U
* device instance $107 r0 *1 -9.5,2 PMOS
M$107 25 20 27 25 PMOS L=1U W=20U AS=40P AD=40P PS=44U PD=44U
* device instance $108 r0 *1 18.5,2 PMOS
M$108 25 20 29 25 PMOS L=1U W=20U AS=40P AD=40P PS=44U PD=44U
* device instance $109 r180 *1 -37.5,-20 HRES
R$109 25 24 1001000 HRES
* device instance $115 m90 *1 75.5,-59.5 D
D$115 35 19 D A=4P P=8U
* device instance $116 r90 *1 63.5,-56 D
D$116 35 20 D A=4P P=8U
* device instance $117 r0 *1 28,-73.5 NMOS
M$117 6 18 19 35 NMOS L=1U W=80U AS=160P AD=160P PS=176U PD=176U
* device instance $121 r0 *1 35,-110.5 NMOS
M$121 9 18 20 35 NMOS L=1U W=80U AS=160P AD=160P PS=176U PD=176U
* device instance $125 r0 *1 -13,-108.5 NMOS
M$125 16 18 18 35 NMOS L=1U W=160U AS=320P AD=320P PS=352U PD=352U
* device instance $133 r0 *1 91.5,-32.5 PMOS
M$133 34 19 18 25 PMOS L=1U W=20U AS=40P AD=40P PS=44U PD=44U
* device instance $134 r0 *1 63.5,-32.5 PMOS
M$134 32 19 18 25 PMOS L=1U W=20U AS=40P AD=40P PS=44U PD=44U
* device instance $135 r0 *1 77.5,-32.5 PMOS
M$135 33 19 18 25 PMOS L=1U W=20U AS=40P AD=40P PS=44U PD=44U
* device instance $136 r0 *1 49.5,-32.5 PMOS
M$136 31 19 18 25 PMOS L=1U W=20U AS=40P AD=40P PS=44U PD=44U
* device instance $137 r0 *1 7.5,-31.5 PMOS
M$137 28 19 20 25 PMOS L=1U W=20U AS=40P AD=40P PS=44U PD=44U
* device instance $138 r0 *1 35.5,-32 PMOS
M$138 30 19 19 25 PMOS L=1U W=20U AS=40P AD=40P PS=44U PD=44U
* device instance $139 r0 *1 21.5,-32 PMOS
M$139 29 20 19 25 PMOS L=1U W=20U AS=40P AD=40P PS=44U PD=44U
* device instance $140 r0 *1 -6.5,-32 PMOS
M$140 27 20 20 25 PMOS L=1U W=20U AS=40P AD=40P PS=44U PD=44U
* device instance $141 r180 *1 -4.5,-212.5 PMOS
M$141 6 6 6 1 PMOS L=1U W=160U AS=320P AD=320P PS=352U PD=352U
* device instance $149 r180 *1 43,-173.5 PMOS
M$149 3 3 3 35 PMOS L=1U W=40U AS=80P AD=80P PS=88U PD=88U
* device instance $151 r180 *1 9.5,-180 PMOS
M$151 9 9 9 5 PMOS L=1U W=20U AS=40P AD=40P PS=44U PD=44U
.ENDS bgr8
