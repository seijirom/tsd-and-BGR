* H:\DESKTOP\ËY¼0SS0\4810\BGR8.ASC
*
*.SUBCKT BGR8 VIN VOUT RES1MEG EXT1MEG R0 R1 R2 R3 VBG
M1 N006 VBG VIN VIN PMOS L=1U W=20U
M2 N004 N001 VIN VIN PMOS L=1U W=20U
M3 N002 N001 VIN VIN PMOS L=1U W=20U
M4 EXT1MEG EXT1MEG VOUT 0 NMOS L=1U W=20U
M5 VBG EXT1MEG N011 0 NMOS L=1U W=20U
M6 N001 EXT1MEG N010 0 NMOS L=1U W=20U
R1 VIN RES1MEG 1MEG
R2 N013 N018 4k
M7 N010 N010 N010 N018 PMOS L=1U W=20U
M8 N011 N011 N011 N013 PMOS L=1U W=20U
M9 N022 N022 N022 0 PMOS L=1U W=20U
M10 N007 VBG VIN VIN PMOS L=1U W=20U
M11 N005 VBG VIN VIN PMOS L=1U W=20U
M12 N003 VBG VIN VIN PMOS L=1U W=20U
M13 N001 N001 N002 VIN PMOS L=1U W=20U
M14 N001 VBG N003 VIN PMOS L=1U W=20U
M15 VBG N001 N004 VIN PMOS L=1U W=20U
M16 VBG VBG N005 VIN PMOS L=1U W=20U
M17 EXT1MEG VBG N006 VIN PMOS L=1U W=20U
M18 EXT1MEG VBG N007 VIN PMOS L=1U W=20U
M19 EXT1MEG EXT1MEG VOUT 0 NMOS L=1U W=20U
M20 EXT1MEG EXT1MEG VOUT 0 NMOS L=1U W=20U
M21 EXT1MEG EXT1MEG VOUT 0 NMOS L=1U W=20U
M22 VBG EXT1MEG N011 0 NMOS L=1U W=20U
M23 VBG EXT1MEG N011 0 NMOS L=1U W=20U
M24 VBG EXT1MEG N011 0 NMOS L=1U W=20U
M25 N001 EXT1MEG N010 0 NMOS L=1U W=20U
M26 N001 EXT1MEG N010 0 NMOS L=1U W=20U
M27 N001 EXT1MEG N010 0 NMOS L=1U W=20U
M28 N011 N011 N011 N013 PMOS L=1U W=20U
M29 N011 N011 N011 N013 PMOS L=1U W=20U
M30 N011 N011 N011 N013 PMOS L=1U W=20U
M31 N011 N011 N011 N013 PMOS L=1U W=20U
M32 N011 N011 N011 N013 PMOS L=1U W=20U
M33 N011 N011 N011 N013 PMOS L=1U W=20U
M34 N011 N011 N011 N013 PMOS L=1U W=20U
R6 0 N023 4k
R7 N019 N023 4k
R8 N019 N024 4k
R9 N020 N024 4k
R10 N020 N025 4k
R11 N021 N025 4k
R12 N021 N018 4k
R4 N012 N014 4k
R14 N014 N015 4k
R15 N015 N016 4k
R16 N016 N017 4k
R17 VOUT R0 4k
R18 VOUT R0 4k
R19 R3 R2 4k
R20 R2 R1 4k
R21 R1 N012 4k
R22 N017 N022 4k
D2 0 N001 D
R3 R3 R2 4k
M35 N022 N022 N022 0 PMOS L=1U W=20U
M36 EXT1MEG EXT1MEG VOUT 0 NMOS L=1U W=20U
M37 EXT1MEG EXT1MEG VOUT 0 NMOS L=1U W=20U
M38 N008 VBG VIN VIN PMOS L=1U W=20U
M39 N009 VBG VIN VIN PMOS L=1U W=20U
M40 EXT1MEG VBG N008 VIN PMOS L=1U W=20U
M41 EXT1MEG VBG N009 VIN PMOS L=1U W=20U
M42 EXT1MEG EXT1MEG VOUT 0 NMOS L=1U W=20U
M43 EXT1MEG EXT1MEG VOUT 0 NMOS L=1U W=20U
R5 0 N023 4k
D1 0 VBG D
*.PARAM RHPO=4K
*.ENDS BGR8

