* Created by KLayout

* cell bgr8
* pin D
* pin R1
* pin Vout
* pin R3
* pin ext1meg
* pin VBG
* pin R2
* pin res1meg
* pin SUBSTRATE
.SUBCKT bgr8 3 4 16 17 18 19 23 24 35
* net 3 D
* net 4 R1
* net 16 Vout
* net 17 R3
* net 18 ext1meg
* net 19 VBG
* net 23 R2
* net 24 res1meg
* net 35 SUBSTRATE
* device instance $3 r0 *1 -45,-108.5 RES
R$3 5 1 4000 RES
* device instance $23 m0 *1 171,-96.5 RES
R$23 23 4 4000 RES
* device instance $53 r0 *1 101,-184.5 RES
R$53 3 4 24000 RES
* device instance $58 m90 *1 -24.5,-199.5 RES
R$58 35 5 26000 RES
* device instance $73 r0 *1 110,-96.5 RES
R$73 16 17 2000 RES
* device instance $83 m90 *1 132,-96.5 RES
R$83 17 23 2000 RES
* device instance $101 r0 *1 88.5,2 PMOS
M$101 25 19 34 25 PMOS L=1U W=20U AS=40P AD=40P PS=44U PD=44U
* device instance $102 r0 *1 74.5,2 PMOS
M$102 25 19 33 25 PMOS L=1U W=20U AS=40P AD=40P PS=44U PD=44U
* device instance $103 r0 *1 32.5,2 PMOS
M$103 25 19 30 25 PMOS L=1U W=20U AS=40P AD=40P PS=44U PD=44U
* device instance $104 r0 *1 60.5,2 PMOS
M$104 25 19 32 25 PMOS L=1U W=20U AS=40P AD=40P PS=44U PD=44U
* device instance $105 r0 *1 46.5,2 PMOS
M$105 25 19 31 25 PMOS L=1U W=20U AS=40P AD=40P PS=44U PD=44U
* device instance $106 r0 *1 4.5,2 PMOS
M$106 25 19 28 25 PMOS L=1U W=20U AS=40P AD=40P PS=44U PD=44U
* device instance $107 r0 *1 -9.5,2 PMOS
M$107 25 20 27 25 PMOS L=1U W=20U AS=40P AD=40P PS=44U PD=44U
* device instance $108 r0 *1 18.5,2 PMOS
M$108 25 20 29 25 PMOS L=1U W=20U AS=40P AD=40P PS=44U PD=44U
* device instance $109 r180 *1 -37.5,-20 HRES
R$109 25 24 1001000 HRES
* device instance $115 m90 *1 75.5,-59.5 D
D$115 35 19 D A=4P P=8U
* device instance $116 r90 *1 63.5,-56 D
D$116 35 20 D A=4P P=8U
* device instance $117 r0 *1 28,-73.5 NMOS
M$117 6 18 19 35 NMOS L=1U W=80U AS=160P AD=160P PS=176U PD=176U
* device instance $121 r0 *1 35,-110.5 NMOS
M$121 9 18 20 35 NMOS L=1U W=80U AS=160P AD=160P PS=176U PD=176U
* device instance $125 r0 *1 -13,-108.5 NMOS
M$125 16 18 18 35 NMOS L=1U W=160U AS=320P AD=320P PS=352U PD=352U
* device instance $133 r0 *1 91.5,-32.5 PMOS
M$133 34 19 18 25 PMOS L=1U W=20U AS=40P AD=40P PS=44U PD=44U
* device instance $134 r0 *1 63.5,-32.5 PMOS
M$134 32 19 18 25 PMOS L=1U W=20U AS=40P AD=40P PS=44U PD=44U
* device instance $135 r0 *1 77.5,-32.5 PMOS
M$135 33 19 18 25 PMOS L=1U W=20U AS=40P AD=40P PS=44U PD=44U
* device instance $136 r0 *1 49.5,-32.5 PMOS
M$136 31 19 18 25 PMOS L=1U W=20U AS=40P AD=40P PS=44U PD=44U
* device instance $137 r0 *1 7.5,-31.5 PMOS
M$137 28 19 20 25 PMOS L=1U W=20U AS=40P AD=40P PS=44U PD=44U
* device instance $138 r0 *1 35.5,-32 PMOS
M$138 30 19 19 25 PMOS L=1U W=20U AS=40P AD=40P PS=44U PD=44U
* device instance $139 r0 *1 21.5,-32 PMOS
M$139 29 20 19 25 PMOS L=1U W=20U AS=40P AD=40P PS=44U PD=44U
* device instance $140 r0 *1 -6.5,-32 PMOS
M$140 27 20 20 25 PMOS L=1U W=20U AS=40P AD=40P PS=44U PD=44U
* device instance $141 r180 *1 -4.5,-212.5 PMOS
M$141 6 6 6 1 PMOS L=1U W=160U AS=320P AD=320P PS=352U PD=352U
* device instance $149 r180 *1 43,-173.5 PMOS
M$149 3 3 3 35 PMOS L=1U W=40U AS=80P AD=80P PS=88U PD=88U
* device instance $151 r180 *1 9.5,-180 PMOS
M$151 9 9 9 5 PMOS L=1U W=20U AS=40P AD=40P PS=44U PD=44U
.ENDS bgr8
