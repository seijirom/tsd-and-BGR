* Created by KLayout

* cell tsd_2021
.SUBCKT tsd_2021
* net 9 SUBSTRATE
* device instance $1 r0 *1 303.5,-218 NMOS
M$1 9 7 4 9 NMOS L=1U W=100U AS=120P AD=120P PS=132U PD=132U
* device instance $6 r0 *1 282.5,-212.5 HRES
R$6 9 3 20000 HRES
* device instance $7 r90 *1 315,-185 HRES
R$7 3 4 100000 HRES
* device instance $10 m90 *1 216.5,-185.5 NMOS
M$10 9 2 1 9 NMOS L=1U W=200U AS=220P AD=220P PS=242U PD=242U
* device instance $20 r0 *1 203.5,-218 NMOS
M$20 9 7 2 9 NMOS L=1U W=200U AS=220P AD=220P PS=242U PD=242U
* device instance $30 r0 *1 252.5,-214 NMOS
M$30 9 21 21 9 NMOS L=1U W=20U AS=40P AD=40P PS=44U PD=44U
* device instance $31 m90 *1 244,-214 NMOS
M$31 9 21 7 9 NMOS L=1U W=20U AS=40P AD=40P PS=44U PD=44U
* device instance $32 r180 *1 266.5,-214 PMOS
M$32 5 5 5 9 PMOS L=1U W=20U AS=40P AD=40P PS=44U PD=44U
* device instance $33 r0 *1 284,-112.5 PMOS
M$33 8 10 14 8 PMOS L=1U W=20U AS=40P AD=40P PS=44U PD=44U
* device instance $34 r180 *1 221,-144 PMOS
M$34 2 10 18 8 PMOS L=1U W=20U AS=40P AD=40P PS=44U PD=44U
* device instance $35 r180 *1 230,-144 PMOS
M$35 2 10 17 8 PMOS L=1U W=20U AS=40P AD=40P PS=44U PD=44U
* device instance $36 r180 *1 243,-143.5 PMOS
M$36 6 10 16 8 PMOS L=1U W=20U AS=40P AD=40P PS=44U PD=44U
* device instance $37 r180 *1 252,-143.5 PMOS
M$37 6 10 15 8 PMOS L=1U W=20U AS=40P AD=40P PS=44U PD=44U
* device instance $38 r180 *1 265,-143.5 PMOS
M$38 5 10 12 8 PMOS L=1U W=20U AS=40P AD=40P PS=44U PD=44U
* device instance $39 r180 *1 274,-143.5 PMOS
M$39 5 10 13 8 PMOS L=1U W=20U AS=40P AD=40P PS=44U PD=44U
* device instance $40 r180 *1 287,-143.5 PMOS
M$40 3 10 14 8 PMOS L=1U W=20U AS=40P AD=40P PS=44U PD=44U
* device instance $41 r180 *1 296,-143.5 PMOS
M$41 3 10 11 8 PMOS L=1U W=20U AS=40P AD=40P PS=44U PD=44U
* device instance $42 r0 *1 218,-113 PMOS
M$42 8 10 18 8 PMOS L=1U W=20U AS=40P AD=40P PS=44U PD=44U
* device instance $43 r0 *1 227,-113 PMOS
M$43 8 10 17 8 PMOS L=1U W=20U AS=40P AD=40P PS=44U PD=44U
* device instance $44 r0 *1 240,-112.5 PMOS
M$44 8 10 16 8 PMOS L=1U W=20U AS=40P AD=40P PS=44U PD=44U
* device instance $45 r0 *1 249,-112.5 PMOS
M$45 8 10 15 8 PMOS L=1U W=20U AS=40P AD=40P PS=44U PD=44U
* device instance $46 r0 *1 262,-112.5 PMOS
M$46 8 10 12 8 PMOS L=1U W=20U AS=40P AD=40P PS=44U PD=44U
* device instance $47 r0 *1 271,-112.5 PMOS
M$47 8 10 13 8 PMOS L=1U W=20U AS=40P AD=40P PS=44U PD=44U
* device instance $48 r0 *1 293,-112.5 PMOS
M$48 8 10 11 8 PMOS L=1U W=20U AS=40P AD=40P PS=44U PD=44U
* device instance $49 m90 *1 253.5,-185 PMOS
M$49 6 5 21 6 PMOS L=1U W=20U AS=40P AD=40P PS=44U PD=44U
* device instance $50 r0 *1 240,-185 PMOS
M$50 6 3 7 6 PMOS L=1U W=20U AS=40P AD=40P PS=44U PD=44U
.ENDS tsd_2021
