* Created by KLayout

* cell bgr_simple
.SUBCKT bgr_simple
* net 1 R1
* net 2 Vdd
* net 8 Vout
* net 9 R0,R3
* net 14 R2
* net 16 SUBSTRATE
* cell instance $2 r0 *1 0,7.5
X$2 15 11 15 12 16 2 2 2 2 2 2 2 2 2 2 2 2 2 2 2 2 2 pch_block
* cell instance $6 r0 *1 -6,-230
X$6 7 16 6 4 13 5 core$BGR
* cell instance $8 r0 *1 -23.5,-92
X$8 15 12 8 11 6 13 16 nch_block
* device instance $1 r0 *1 176.5,-184.5 RES
R$1 97 54 800
* device instance $2 r0 *1 172.5,-184.5 RES
R$2 97 55 800
* device instance $3 r0 *1 168.5,-184.5 RES
R$3 99 55 800
* device instance $4 r0 *1 164.5,-184.5 RES
R$4 99 43 800
* device instance $5 r0 *1 160.5,-184.5 RES
R$5 88 43 800
* device instance $6 r0 *1 157,-184.5 RES
R$6 88 44 800
* device instance $7 r0 *1 153,-184.5 RES
R$7 89 44 800
* device instance $8 r0 *1 149,-184.5 RES
R$8 89 45 800
* device instance $9 r0 *1 145,-184.5 RES
R$9 90 45 800
* device instance $10 r0 *1 141,-184.5 RES
R$10 90 46 800
* device instance $11 r0 *1 137.5,-184.5 RES
R$11 91 46 800
* device instance $12 r0 *1 133.5,-184.5 RES
R$12 91 47 800
* device instance $13 r0 *1 129.5,-184.5 RES
R$13 92 47 800
* device instance $14 r0 *1 125.5,-184.5 RES
R$14 92 48 800
* device instance $15 r0 *1 121.5,-184.5 RES
R$15 98 48 800
* device instance $16 r0 *1 118,-184.5 RES
R$16 98 50 800
* device instance $17 r0 *1 114,-184.5 RES
R$17 93 50 800
* device instance $18 r0 *1 110,-184.5 RES
R$18 93 51 800
* device instance $19 r0 *1 106,-184.5 RES
R$19 94 51 800
* device instance $20 r0 *1 102,-184.5 RES
R$20 94 52 800
* device instance $21 r0 *1 98,-184.5 RES
R$21 95 52 800
* device instance $22 r0 *1 94,-184.5 RES
R$22 95 53 800
* device instance $23 r0 *1 82,-184.5 RES
R$23 7 20 800
* device instance $24 r0 *1 86,-184.5 RES
R$24 96 20 800
* device instance $25 r0 *1 90,-184.5 RES
R$25 96 53 800
* device instance $26 r0 *1 -131,-175.5 RES
R$26 101 57 800
* device instance $27 r0 *1 -127,-175.5 RES
R$27 101 58 800
* device instance $28 r0 *1 -123,-175.5 RES
R$28 102 58 800
* device instance $29 r0 *1 -119,-175.5 RES
R$29 102 59 800
* device instance $30 r0 *1 -115,-175.5 RES
R$30 103 59 800
* device instance $31 r0 *1 -111,-175.5 RES
R$31 103 60 800
* device instance $32 r0 *1 -107,-175.5 RES
R$32 109 60 800
* device instance $33 r0 *1 -103,-175.5 RES
R$33 109 66 800
* device instance $34 r0 *1 -99,-175.5 RES
R$34 108 66 800
* device instance $35 r0 *1 -95,-175.5 RES
R$35 108 65 800
* device instance $36 r0 *1 -91,-175.5 RES
R$36 107 65 800
* device instance $37 r0 *1 -87,-175.5 RES
R$37 107 64 800
* device instance $38 r0 *1 -83,-175.5 RES
R$38 106 64 800
* device instance $39 r0 *1 -79,-175.5 RES
R$39 106 63 800
* device instance $40 r0 *1 -75,-175.5 RES
R$40 16 63 800
* device instance $41 r0 *1 -71,-175.5 RES
R$41 105 65 800
* device instance $42 r0 *1 -67,-175.5 RES
R$42 105 62 800
* device instance $43 r0 *1 -63,-175.5 RES
R$43 104 62 800
* device instance $44 r0 *1 -59,-175.5 RES
R$44 104 49 800
* device instance $45 r0 *1 -55,-175.5 RES
R$45 16 49 800
* device instance $46 r0 *1 201.5,-97.5 RES
R$46 77 1 800
* device instance $47 r0 *1 197.5,-97.5 RES
R$47 77 33 800
* device instance $48 r0 *1 193.5,-97.5 RES
R$48 78 33 800
* device instance $49 r0 *1 189.5,-97.5 RES
R$49 78 34 800
* device instance $50 r0 *1 185.5,-97.5 RES
R$50 54 34 800
* device instance $51 r0 *1 179,-96.5 RES
R$51 1 22 800
* device instance $52 r0 *1 82,-96.5 RES
R$52 8 35 800
* device instance $53 r0 *1 86,-96.5 RES
R$53 79 35 800
* device instance $54 r0 *1 90,-96.5 RES
R$54 79 36 800
* device instance $55 r0 *1 94,-96.5 RES
R$55 80 36 800
* device instance $56 r0 *1 98,-96.5 RES
R$56 80 9 800
* device instance $57 r0 *1 102,-96.5 RES
R$57 8 37 800
* device instance $58 r0 *1 106,-96.5 RES
R$58 87 37 800
* device instance $59 r0 *1 110,-96.5 RES
R$59 87 38 800
* device instance $60 r0 *1 114,-96.5 RES
R$60 82 38 800
* device instance $61 r0 *1 118,-96.5 RES
R$61 82 9 800
* device instance $62 r0 *1 124,-96.5 RES
R$62 83 14 800
* device instance $63 r0 *1 128,-96.5 RES
R$63 83 39 800
* device instance $64 r0 *1 132,-96.5 RES
R$64 84 39 800
* device instance $65 r0 *1 136,-96.5 RES
R$65 84 40 800
* device instance $66 r0 *1 140,-96.5 RES
R$66 9 40 800
* device instance $67 r0 *1 143.5,-96.5 RES
R$67 9 41 800
* device instance $68 r0 *1 147.5,-96.5 RES
R$68 85 41 800
* device instance $69 r0 *1 151.5,-96.5 RES
R$69 85 42 800
* device instance $70 r0 *1 155.5,-96.5 RES
R$70 86 42 800
* device instance $71 r0 *1 159.5,-96.5 RES
R$71 86 14 800
* device instance $72 r0 *1 163,-96.5 RES
R$72 81 14 800
* device instance $73 r0 *1 167,-96.5 RES
R$73 81 21 800
* device instance $74 r0 *1 171,-96.5 RES
R$74 67 21 800
* device instance $75 r0 *1 175,-96.5 RES
R$75 67 22 800
* device instance $76 r0 *1 -131,-87.5 RES
R$76 57 23 800
* device instance $77 r0 *1 -127,-87.5 RES
R$77 68 23 800
* device instance $78 r0 *1 -123,-87.5 RES
R$78 68 24 800
* device instance $79 r0 *1 -119,-87.5 RES
R$79 69 24 800
* device instance $80 r0 *1 -115,-87.5 RES
R$80 69 25 800
* device instance $81 r0 *1 -111,-87.5 RES
R$81 70 25 800
* device instance $82 r0 *1 -107,-87.5 RES
R$82 70 26 800
* device instance $83 r0 *1 -103,-87.5 RES
R$83 71 26 800
* device instance $84 r0 *1 -99,-87.5 RES
R$84 71 27 800
* device instance $85 r0 *1 -95,-87.5 RES
R$85 76 27 800
* device instance $86 r0 *1 -91,-87.5 RES
R$86 76 28 800
* device instance $87 r0 *1 -87,-87.5 RES
R$87 72 28 800
* device instance $88 r0 *1 -83,-87.5 RES
R$88 72 29 800
* device instance $89 r0 *1 -79,-87.5 RES
R$89 73 29 800
* device instance $90 r0 *1 -75,-87.5 RES
R$90 73 30 800
* device instance $91 r0 *1 -71,-87.5 RES
R$91 74 30 800
* device instance $92 r0 *1 -67,-87.5 RES
R$92 74 31 800
* device instance $93 r0 *1 -63,-87.5 RES
R$93 75 31 800
* device instance $94 r0 *1 -59,-87.5 RES
R$94 75 32 800
* device instance $95 r0 *1 -55,-87.5 RES
R$95 4 32 800
* device instance $96 r0 *1 -51.5,-87.5 RES
R$96 4 61 800
* device instance $97 r0 *1 -47.5,-87.5 RES
R$97 100 61 800
* device instance $98 r0 *1 -43.5,-87.5 RES
R$98 100 56 800
* device instance $99 r0 *1 -39.5,-87.5 RES
R$99 3 56 800
* device instance $100 r0 *1 -35.5,-87.5 RES
R$100 3 5 800
* device instance $101 r0 *1 -52.5,15.5 HRES
R$101 19 10 245000
* device instance $102 r0 *1 -48.5,16.5 HRES
R$102 19 17 252000
* device instance $103 r0 *1 -44.5,16.5 HRES
R$103 18 17 252000
* device instance $104 r0 *1 -40.5,16.5 HRES
R$104 18 2 252000
.ENDS bgr_simple

* cell nch_block
* pin 
* pin 
* pin 
* pin 
* pin 
* pin 
* pin SUBSTRATE
.SUBCKT nch_block 1 2 3 4 5 6 7
* net 7 SUBSTRATE
* cell instance $1 r0 *1 56,-1
X$1 5 1 2 7 Nch
* cell instance $2 r0 *1 24.5,34.5
X$2 5 1 2 7 Nch
* cell instance $3 r0 *1 37,34
X$3 5 1 2 7 Nch
* cell instance $4 r0 *1 68,-1
X$4 5 1 2 7 Nch
* cell instance $8 r0 *1 8,-1
X$8 3 2 2 7 Nch
* cell instance $9 r0 *1 49,34
X$9 6 4 2 7 Nch
* cell instance $10 r0 *1 1,34
X$10 3 2 2 7 Nch
* cell instance $11 r0 *1 13,34
X$11 3 2 2 7 Nch
* cell instance $12 r0 *1 61,34
X$12 6 4 2 7 Nch
* cell instance $13 r0 *1 85,34
X$13 3 2 2 7 Nch
* cell instance $14 r0 *1 73,34
X$14 3 2 2 7 Nch
* cell instance $15 r0 *1 92,-1
X$15 3 2 2 7 Nch
* cell instance $16 r0 *1 80,-1
X$16 3 2 2 7 Nch
* cell instance $17 r0 *1 32,-1
X$17 6 4 2 7 Nch
* cell instance $18 r0 *1 44,-1
X$18 6 4 2 7 Nch
* cell instance $19 r0 *1 20,-1
X$19 3 2 2 7 Nch
.ENDS nch_block

* cell pch_block
* pin 
* pin 
* pin 
* pin 
* pin 
* pin 
* pin 
* pin 
* pin 
* pin 
* pin 
* pin 
* pin 
* pin 
* pin 
* pin 
* pin 
* pin 
* pin 
* pin 
* pin 
* pin 
.SUBCKT pch_block 1 2 3 4 5 6 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30
* cell instance $1 r0 *1 1,-44.5
X$1 1 5 protection$1
* cell instance $3 r0 *1 -12,30
X$3 30 13 1 22 Pch
* cell instance $4 r0 *1 -9,-4
X$4 13 1 1 6 Pch
* cell instance $5 r0 *1 5,-3.5
X$5 8 1 2 6 Pch
* cell instance $6 r0 *1 93,-38
X$6 2 5 protection
* cell instance $14 r0 *1 86,30
X$14 24 10 2 16 Pch
* cell instance $15 r0 *1 61,-4.5
X$15 12 4 2 6 Pch
* cell instance $16 r0 *1 47,-4.5
X$16 14 4 2 6 Pch
* cell instance $17 r0 *1 33,-4.5
X$17 7 2 2 6 Pch
* cell instance $18 r0 *1 2,30
X$18 25 8 2 17 Pch
* cell instance $19 r0 *1 44,30
X$19 26 14 2 18 Pch
* cell instance $20 r0 *1 58,30
X$20 27 12 2 19 Pch
* cell instance $21 r0 *1 30,30
X$21 28 7 2 20 Pch
* cell instance $22 r0 *1 72,30
X$22 29 11 2 21 Pch
* cell instance $23 r0 *1 75,-4.5
X$23 11 4 2 6 Pch
* cell instance $24 r0 *1 89,-4.5
X$24 10 4 2 6 Pch
* cell instance $25 r0 *1 19,-4
X$25 9 2 3 6 Pch
* cell instance $27 r0 *1 16,30
X$27 23 9 3 15 Pch
.ENDS pch_block

* cell core$BGR
* pin 
* pin 
* pin 
* pin 
* pin 
* pin 
.SUBCKT core$BGR 1 2 3 4 5 6
* cell instance $1 r180 *1 54.5,38.5
X$1 1 2 pchdiode
* cell instance $2 r180 *1 54.5,73
X$2 1 2 pchdiode
* cell instance $3 r180 *1 32.5,50.5
X$3 6 5 3 4 diodeblock
.ENDS core$BGR

* cell Nch
* pin 
* pin 
* pin 
* pin SUBSTRATE
.SUBCKT Nch 1 2 3 4
* net 4 SUBSTRATE
* device instance $1 r0 *1 2.5,13 NMOS
M$1 1 3 2 4 NMOS L=1U W=20U AS=40P AD=40P PS=44U PD=44U
.ENDS Nch

* cell protection
* pin 
* pin 
.SUBCKT protection 1 2
* device instance $1 r0 *1 4.5,24 D
D$1 2 1 D A=1P P=4U
.ENDS protection

* cell protection$1
* pin 
* pin 
.SUBCKT protection$1 1 2
* device instance $1 r0 *1 4,24 D
D$1 2 1 D A=1P P=4U
.ENDS protection$1

* cell diodeblock
* pin 
* pin 
* pin 
* pin 
.SUBCKT diodeblock 1 2 3 4
* cell instance $1 r0 *1 -2.5,-33.5
X$1 2 1 pchdiode
* cell instance $2 r0 *1 25.5,-71
X$2 2 1 pchdiode
* cell instance $3 r0 *1 11,-71
X$3 2 1 pchdiode
* cell instance $4 r0 *1 -2.5,-71
X$4 2 1 pchdiode
* cell instance $5 r0 *1 25.5,-33.5
X$5 2 1 pchdiode
* cell instance $6 r0 *1 25.5,4
X$6 2 1 pchdiode
* cell instance $7 r0 *1 11,4
X$7 2 1 pchdiode
* cell instance $8 r0 *1 -2.5,4
X$8 2 1 pchdiode
* cell instance $9 r0 *1 11,-33.5
X$9 3 4 pchdiode
.ENDS diodeblock

* cell pchdiode
* pin 
* pin 
.SUBCKT pchdiode 1 2
* cell instance $1 r0 *1 2,1
X$1 2 1 1 1 pch1x20
.ENDS pchdiode

* cell pch1x20
* pin 
* pin 
* pin 
* pin 
.SUBCKT pch1x20 1 2 3 4
* cell instance $1 r0 *1 1,2.5
X$1 4 3 2 1 Pch
.ENDS pch1x20

* cell Pch
* pin 
* pin 
* pin 
* pin 
.SUBCKT Pch 1 2 3 4
* device instance $1 r0 *1 2.5,13 PMOS
M$1 1 3 2 4 PMOS L=1U W=20U AS=40P AD=40P PS=44U PD=44U
.ENDS Pch
