* Created by KLayout

* cell bgr_simple
.SUBCKT bgr_simple
* net 1 Vout
* net 2 Vin
* net 5 R2
* net 6 R1
* net 11 D
* net 12 R3
* net 26 Gnd
* cell instance $3 r0 *1 12,-43
X$3 2 8 10 2 pch1x20
* cell instance $4 r0 *1 3,-43
X$4 2 8 8 2 pch1x20
* cell instance $5 r0 *1 21,-43
X$5 2 10 7 2 pch1x20
* cell instance $6 r0 *1 30,-43
X$6 2 10 7 2 pch1x20
* cell instance $7 r180 *1 39.5,-151.5
X$7 13 25 9 3 diodeblock
* cell instance $8 r0 *1 3,-78
X$8 26 7 3 8 nch1x20
* cell instance $9 r0 *1 21,-78
X$9 26 7 4 7 nch1x20
* cell instance $10 r0 *1 30,-78
X$10 26 7 4 7 nch1x20
* cell instance $16 r0 *1 12,-78
X$16 26 7 13 10 nch1x20
* cell instance $17 r270 *1 3,-43
X$17 26 protection
* cell instance $18 r90 *1 26.5,-53
X$18 26 protection
* cell instance $21 m45 *1 -11.5,-53
X$21 26 protection
* cell instance $23 r180 *1 57.5,-157.5
X$23 11 26 pchdiode
* cell instance $24 r180 *1 57.5,-123
X$24 11 26 pchdiode
* device instance $1 r0 *1 -87.5,-147.5 RES
R$1 69 22 800
* device instance $2 r0 *1 -83.5,-147.5 RES
R$2 69 44 800
* device instance $3 r0 *1 -79.5,-147.5 RES
R$3 84 44 800
* device instance $4 r0 *1 -75.5,-147.5 RES
R$4 84 45 800
* device instance $5 r0 *1 -71.5,-147.5 RES
R$5 23 45 800
* device instance $6 r0 *1 -67.5,-147.5 RES
R$6 23 46 800
* device instance $7 r0 *1 -63.5,-147.5 RES
R$7 85 46 800
* device instance $8 r0 *1 -59.5,-147.5 RES
R$8 85 47 800
* device instance $9 r0 *1 -55.5,-147.5 RES
R$9 86 47 800
* device instance $10 r0 *1 -51.5,-147.5 RES
R$10 86 24 800
* device instance $11 r0 *1 -47.5,-147.5 RES
R$11 91 24 800
* device instance $12 r0 *1 -43.5,-147.5 RES
R$12 91 49 800
* device instance $13 r0 *1 -39.5,-147.5 RES
R$13 87 49 800
* device instance $14 r0 *1 -35.5,-147.5 RES
R$14 87 50 800
* device instance $15 r0 *1 -31.5,-147.5 RES
R$15 26 50 800
* device instance $16 r0 *1 -27.5,-147.5 RES
R$16 88 9 800
* device instance $17 r0 *1 -23.5,-147.5 RES
R$17 88 51 800
* device instance $18 r0 *1 -19.5,-147.5 RES
R$18 89 51 800
* device instance $19 r0 *1 -15.5,-147.5 RES
R$19 89 52 800
* device instance $20 r0 *1 -11.5,-147.5 RES
R$20 25 52 800
* device instance $21 r0 *1 166.5,-147.5 RES
R$21 90 12 800
* device instance $22 r0 *1 162.5,-147.5 RES
R$22 90 40 800
* device instance $23 r0 *1 158.5,-147.5 RES
R$23 83 40 800
* device instance $24 r0 *1 154.5,-147.5 RES
R$24 83 39 800
* device instance $25 r0 *1 150.5,-147.5 RES
R$25 18 39 800
* device instance $26 r0 *1 146.5,-147.5 RES
R$26 18 38 800
* device instance $27 r0 *1 142.5,-147.5 RES
R$27 77 38 800
* device instance $28 r0 *1 138.5,-147.5 RES
R$28 77 48 800
* device instance $29 r0 *1 70.5,-147.5 RES
R$29 11 37 800
* device instance $30 r0 *1 74.5,-147.5 RES
R$30 76 37 800
* device instance $31 r0 *1 78.5,-147.5 RES
R$31 76 36 800
* device instance $32 r0 *1 82.5,-147.5 RES
R$32 75 36 800
* device instance $33 r0 *1 86.5,-147.5 RES
R$33 75 15 800
* device instance $34 r0 *1 90.5,-147.5 RES
R$34 78 15 800
* device instance $35 r0 *1 94.5,-147.5 RES
R$35 78 35 800
* device instance $36 r0 *1 98.5,-147.5 RES
R$36 79 35 800
* device instance $37 r0 *1 102.5,-147.5 RES
R$37 79 41 800
* device instance $38 r0 *1 106.5,-147.5 RES
R$38 16 41 800
* device instance $39 r0 *1 110.5,-147.5 RES
R$39 16 42 800
* device instance $40 r0 *1 114.5,-147.5 RES
R$40 80 42 800
* device instance $41 r0 *1 118.5,-147.5 RES
R$41 80 43 800
* device instance $42 r0 *1 122.5,-147.5 RES
R$42 81 43 800
* device instance $43 r0 *1 126.5,-147.5 RES
R$43 81 17 800
* device instance $44 r0 *1 130.5,-147.5 RES
R$44 82 17 800
* device instance $45 r0 *1 134.5,-147.5 RES
R$45 82 48 800
* device instance $46 r0 *1 -87.5,-59.5 RES
R$46 22 73 800
* device instance $47 r0 *1 -83.5,-59.5 RES
R$47 99 73 800
* device instance $48 r0 *1 -79.5,-59.5 RES
R$48 99 62 800
* device instance $49 r0 *1 -75.5,-59.5 RES
R$49 100 62 800
* device instance $50 r0 *1 -71.5,-59.5 RES
R$50 100 14 800
* device instance $51 r0 *1 -67.5,-59.5 RES
R$51 34 14 800
* device instance $52 r0 *1 -63.5,-59.5 RES
R$52 34 63 800
* device instance $53 r0 *1 -59.5,-59.5 RES
R$53 101 63 800
* device instance $54 r0 *1 -55.5,-59.5 RES
R$54 101 64 800
* device instance $55 r0 *1 -51.5,-59.5 RES
R$55 21 64 800
* device instance $56 r0 *1 -47.5,-59.5 RES
R$56 21 74 800
* device instance $57 r0 *1 -43.5,-59.5 RES
R$57 102 74 800
* device instance $58 r0 *1 -39.5,-59.5 RES
R$58 102 68 800
* device instance $59 r0 *1 -35.5,-59.5 RES
R$59 105 68 800
* device instance $60 r0 *1 -31.5,-59.5 RES
R$60 105 20 800
* device instance $61 r0 *1 -27.5,-59.5 RES
R$61 104 20 800
* device instance $62 r0 *1 -23.5,-59.5 RES
R$62 104 66 800
* device instance $63 r0 *1 -19.5,-59.5 RES
R$63 103 66 800
* device instance $64 r0 *1 -15.5,-59.5 RES
R$64 103 65 800
* device instance $65 r0 *1 -11.5,-59.5 RES
R$65 19 65 800
* device instance $66 r0 *1 -7.5,-59.5 RES
R$66 19 9 800
* device instance $67 r0 *1 166.5,-59.5 RES
R$67 12 67 800
* device instance $68 r0 *1 162.5,-59.5 RES
R$68 95 67 800
* device instance $69 r0 *1 158.5,-59.5 RES
R$69 95 53 800
* device instance $70 r0 *1 154.5,-59.5 RES
R$70 70 53 800
* device instance $71 r0 *1 150.5,-59.5 RES
R$71 70 5 800
* device instance $72 r0 *1 146.5,-59.5 RES
R$72 92 5 800
* device instance $73 r0 *1 142.5,-59.5 RES
R$73 92 54 800
* device instance $74 r0 *1 138.5,-59.5 RES
R$74 98 54 800
* device instance $75 r0 *1 70.5,-59.5 RES
R$75 6 55 800
* device instance $76 r0 *1 74.5,-59.5 RES
R$76 93 55 800
* device instance $77 r0 *1 78.5,-59.5 RES
R$77 93 56 800
* device instance $78 r0 *1 82.5,-59.5 RES
R$78 94 56 800
* device instance $79 r0 *1 86.5,-59.5 RES
R$79 94 4 800
* device instance $80 r0 *1 90.5,-59.5 RES
R$80 72 4 800
* device instance $81 r0 *1 94.5,-59.5 RES
R$81 72 57 800
* device instance $82 r0 *1 98.5,-59.5 RES
R$82 96 57 800
* device instance $83 r0 *1 102.5,-59.5 RES
R$83 96 58 800
* device instance $84 r0 *1 106.5,-59.5 RES
R$84 6 58 800
* device instance $85 r0 *1 110.5,-59.5 RES
R$85 71 5 800
* device instance $86 r0 *1 114.5,-59.5 RES
R$86 71 59 800
* device instance $87 r0 *1 118.5,-59.5 RES
R$87 97 59 800
* device instance $88 r0 *1 122.5,-59.5 RES
R$88 97 60 800
* device instance $89 r0 *1 126.5,-59.5 RES
R$89 6 60 800
* device instance $90 r0 *1 130.5,-59.5 RES
R$90 6 61 800
* device instance $91 r0 *1 134.5,-59.5 RES
R$91 98 61 800
* device instance $92 r0 *1 64.5,-21.5 RES
R$92 28 4 200
* device instance $93 r0 *1 60.5,-21.5 RES
R$93 28 30 200
* device instance $94 r0 *1 56.5,-21.5 RES
R$94 27 30 200
* device instance $95 r0 *1 52.5,-21.5 RES
R$95 27 29 200
* device instance $96 r0 *1 48.5,-21.5 RES
R$96 1 29 200
* device instance $97 r0 *1 59.5,-80 HRES
R$97 33 2 262500
* device instance $98 r0 *1 55.5,-80 HRES
R$98 33 31 262500
* device instance $99 r0 *1 51.5,-80 HRES
R$99 32 31 262500
* device instance $100 r0 *1 47.5,-80 HRES
R$100 32 7 262500
.ENDS bgr_simple

* cell protection
* pin 
.SUBCKT protection 2
* device instance $1 r0 *1 4.5,24 D
D$1 2 1 D A=1P P=4U
.ENDS protection

* cell diodeblock
* pin 
* pin 
* pin 
* pin 
.SUBCKT diodeblock 1 2 3 4
* cell instance $1 r0 *1 -2.5,-71
X$1 1 2 pchdiode
* cell instance $2 r0 *1 25.5,-71
X$2 1 2 pchdiode
* cell instance $3 r0 *1 11,-71
X$3 1 2 pchdiode
* cell instance $4 r0 *1 25.5,-33.5
X$4 1 2 pchdiode
* cell instance $5 r0 *1 -2.5,-33.5
X$5 1 2 pchdiode
* cell instance $6 r0 *1 25.5,4
X$6 1 2 pchdiode
* cell instance $7 r0 *1 11,4
X$7 1 2 pchdiode
* cell instance $8 r0 *1 -2.5,4
X$8 1 2 pchdiode
* cell instance $9 r0 *1 11,-33.5
X$9 4 3 pchdiode
.ENDS diodeblock

* cell nch1x20
* pin SUBSTRATE
* pin 
* pin 
* pin 
.SUBCKT nch1x20 1 2 3 4
* net 1 SUBSTRATE
* cell instance $1 r0 *1 0.5,-0.5
X$1 3 4 2 1 Nch
.ENDS nch1x20

* cell Nch
* pin 
* pin 
* pin 
* pin SUBSTRATE
.SUBCKT Nch 1 2 3 4
* net 4 SUBSTRATE
* device instance $1 r0 *1 2.5,13 NMOS
M$1 1 3 2 4 NMOS L=1U W=20U AS=40P AD=40P PS=44U PD=44U
.ENDS Nch

* cell pchdiode
* pin 
* pin 
.SUBCKT pchdiode 1 2
* cell instance $1 r0 *1 2,1
X$1 2 1 1 1 pch1x20
.ENDS pchdiode

* cell pch1x20
* pin 
* pin 
* pin 
* pin 
.SUBCKT pch1x20 1 2 3 4
* cell instance $1 r0 *1 1,2.5
X$1 4 3 2 1 Pch
.ENDS pch1x20

* cell Pch
* pin 
* pin 
* pin 
* pin 
.SUBCKT Pch 1 2 3 4
* device instance $1 r0 *1 2.5,13 PMOS
M$1 1 3 2 4 PMOS L=1U W=20U AS=40P AD=40P PS=44U PD=44U
.ENDS Pch
