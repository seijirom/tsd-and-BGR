* Z:\HOME\SEIJIROM\WORK\2021_9\TSD_AND_BGR\TSD_TB_WITH_RESISTORS.ASC
*XX2 N003 N004 N002 NC_01 N012 N009 N008 N005 N007 BGR8
*V1 N001 0 5
R1 N011 NC_02 25K
R2 N011 NC_03 35K
R3 N011 NC_04 50K
R4 N011 NC_05 65K
R5 N011 NC_06 75K
*V2 N003 0 5
XX1 N001 N007 NC_07 N011 N010 N006 N006 0 TSD_CORE
*
* BLOCK SYMBOL DEFINITIONS
.SUBCKT BGR8 VIN VOUT RES1MEG EXT1MEG D R1 R2 R3 VBG
M19 N006 VBG VIN VIN PMOS L=1U W=20U
M17 N004 N001 VIN VIN PMOS L=1U W=20U
M11 N002 N001 VIN VIN PMOS L=1U W=20U
M35 EXT1MEG EXT1MEG VOUT 0 NMOS L=1U W=20U
M31 VBG EXT1MEG N011 0 NMOS L=1U W=20U
M27 N001 EXT1MEG N010 0 NMOS L=1U W=20U
R1 VIN RES1MEG 1MEG
R2 N013 N018 4K
M47 N010 N010 N010 N018 PMOS L=1U W=20U
M45 N011 N011 N011 N013 PMOS L=1U W=20U
M53 D D D 0 PMOS L=1U W=20U
M22 N007 VBG VIN VIN PMOS L=1U W=20U
M18 N005 VBG VIN VIN PMOS L=1U W=20U
M12 N003 VBG VIN VIN PMOS L=1U W=20U
M13 N001 N001 N002 VIN PMOS L=1U W=20U
M14 N001 VBG N003 VIN PMOS L=1U W=20U
M15 VBG N001 N004 VIN PMOS L=1U W=20U
M16 VBG VBG N005 VIN PMOS L=1U W=20U
M20 EXT1MEG VBG N006 VIN PMOS L=1U W=20U
M21 EXT1MEG VBG N007 VIN PMOS L=1U W=20U
M36 EXT1MEG EXT1MEG VOUT 0 NMOS L=1U W=20U
M23 EXT1MEG EXT1MEG VOUT 0 NMOS L=1U W=20U
M24 EXT1MEG EXT1MEG VOUT 0 NMOS L=1U W=20U
M32 VBG EXT1MEG N011 0 NMOS L=1U W=20U
M28 VBG EXT1MEG N011 0 NMOS L=1U W=20U
M29 VBG EXT1MEG N011 0 NMOS L=1U W=20U
M30 N001 EXT1MEG N010 0 NMOS L=1U W=20U
M33 N001 EXT1MEG N010 0 NMOS L=1U W=20U
M34 N001 EXT1MEG N010 0 NMOS L=1U W=20U
M43 N011 N011 N011 N013 PMOS L=1U W=20U
M46 N011 N011 N011 N013 PMOS L=1U W=20U
M49 N011 N011 N011 N013 PMOS L=1U W=20U
M48 N011 N011 N011 N013 PMOS L=1U W=20U
M50 N011 N011 N011 N013 PMOS L=1U W=20U
M44 N011 N011 N011 N013 PMOS L=1U W=20U
M51 N011 N011 N011 N013 PMOS L=1U W=20U
R6 0 N022 4K
R7 N019 N022 4K
R8 N019 N023 4K
R9 N020 N023 4K
R10 N020 N024 4K
R11 N021 N024 4K
R12 N021 N018 4K
R4 N012 N014 4K
R14 N014 N015 4K
R15 N015 N016 4K
R16 N016 N017 4K
R17 VOUT R3 4K
R18 VOUT R3 4K
R19 R3 R2 4K
R20 R2 R1 4K
R21 R1 N012 4K
R22 N017 D 4K
D2 0 N001 D
R3 R3 R2 4K
M52 D D D 0 PMOS L=1U W=20U
M37 EXT1MEG EXT1MEG VOUT 0 NMOS L=1U W=20U
M38 EXT1MEG EXT1MEG VOUT 0 NMOS L=1U W=20U
M42 N008 VBG VIN VIN PMOS L=1U W=20U
M39 N009 VBG VIN VIN PMOS L=1U W=20U
M40 EXT1MEG VBG N008 VIN PMOS L=1U W=20U
M41 EXT1MEG VBG N009 VIN PMOS L=1U W=20U
M25 EXT1MEG EXT1MEG VOUT 0 NMOS L=1U W=20U
M26 EXT1MEG EXT1MEG VOUT 0 NMOS L=1U W=20U
R5 0 N022 4K
D1 0 VBG D
*.PARAM RHPO=4K
.ENDS BGR8
*
.SUBCKT TSD_CORE VIN VBGR TSD A B C R100K R20K
M23 A VBGR N008 VIN PMOS L=1U W=20U
R6 A R20K 20K
M29 B VBGR N005 VIN PMOS L=1U W=20U
M12 B B B 0 PMOS L=1U W=20U
M33 N009 VBGR N003 VIN PMOS L=1U W=20U
M14 N012 B N009 N009 PMOS L=1U W=20U
M15 N011 A N009 N009 PMOS L=1U W=20U
M16 N011 N012 0 0 NMOS L=1U W=20U
M17 N012 N012 0 0 NMOS L=1U W=20U
M21 C N011 0 0 NMOS L=1U W=100U
M22 N008 VBGR VIN VIN PMOS L=1U W=20U
M28 N005 VBGR VIN VIN PMOS L=1U W=20U
M32 N003 VBGR VIN VIN PMOS L=1U W=20U
M31 N009 VBGR N004 VIN PMOS L=1U W=20U
M30 N004 VBGR VIN VIN PMOS L=1U W=20U
M27 B VBGR N006 VIN PMOS L=1U W=20U
M26 N006 VBGR VIN VIN PMOS L=1U W=20U
M25 A VBGR N007 VIN PMOS L=1U W=20U
M24 N007 VBGR VIN VIN PMOS L=1U W=20U
R7 A R100K 100K
M19 N010 N011 0 0 NMOS L=1U W=200U
M1 N010 VBGR N001 VIN PMOS L=1U W=20U
M2 N001 VBGR VIN VIN PMOS L=1U W=20U
M3 N010 VBGR N002 VIN PMOS L=1U W=20U
M4 N002 VBGR VIN VIN PMOS L=1U W=20U
M5 TSD N010 0 0 NMOS L=1U W=200U
*.INCLUDE "./MODELS/OR1_MOS"
.ENDS TSD_CORE

.MODEL D D
.LIB C:\USERS\SEIJIROM\MY DOCUMENTS\LTSPICEXVII\LIB\CMP\STANDARD.DIO
.MODEL NMOS NMOS
.MODEL PMOS PMOS
.LIB C:\USERS\SEIJIROM\MY DOCUMENTS\LTSPICEXVII\LIB\CMP\STANDARD.MOS
* D*2: A=1 B=28K
* D*3:A=1 B=42K
.DC TEMP _50 150 0.1
*.INCLUDE "./MODELS/OR1_MOS"
;STEP PARAM VDD 3.5 5 0.5
.BACKANNO
.GLOBAL 0
.END
