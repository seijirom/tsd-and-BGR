* Created by KLayout

* cell tsd_2021
.SUBCKT tsd_2021
* net 9 SUBSTRATE
* device instance $1 r0 *1 186,-218 NMOS
M$1 9 7 3 9 NMOS L=1U W=200U AS=220P AD=220P PS=242U PD=242U
* device instance $11 r0 *1 286,-218 NMOS
M$11 9 7 4 9 NMOS L=1U W=100U AS=120P AD=120P PS=132U PD=132U
* device instance $16 r0 *1 266,-202.5 HRES
R$16 9 1 20000 HRES
* device instance $17 r90 *1 297.5,-185 HRES
R$17 1 4 100000 HRES
* device instance $20 m90 *1 206.5,-185.5 NMOS
M$20 9 3 2 9 NMOS L=1U W=200U AS=220P AD=220P PS=242U PD=242U
* device instance $30 r0 *1 266.5,-112.5 PMOS
M$30 8 10 14 8 PMOS L=1U W=20U AS=40P AD=40P PS=44U PD=44U
* device instance $31 r0 *1 200.5,-112.5 PMOS
M$31 8 10 18 8 PMOS L=1U W=20U AS=40P AD=40P PS=44U PD=44U
* device instance $32 r0 *1 209.5,-112.5 PMOS
M$32 8 10 17 8 PMOS L=1U W=20U AS=40P AD=40P PS=44U PD=44U
* device instance $33 r0 *1 222.5,-112.5 PMOS
M$33 8 10 16 8 PMOS L=1U W=20U AS=40P AD=40P PS=44U PD=44U
* device instance $34 r0 *1 231.5,-112.5 PMOS
M$34 8 10 15 8 PMOS L=1U W=20U AS=40P AD=40P PS=44U PD=44U
* device instance $35 r0 *1 244.5,-112.5 PMOS
M$35 8 10 12 8 PMOS L=1U W=20U AS=40P AD=40P PS=44U PD=44U
* device instance $36 r0 *1 253.5,-112.5 PMOS
M$36 8 10 13 8 PMOS L=1U W=20U AS=40P AD=40P PS=44U PD=44U
* device instance $37 r0 *1 275.5,-112.5 PMOS
M$37 8 10 11 8 PMOS L=1U W=20U AS=40P AD=40P PS=44U PD=44U
* device instance $38 r0 *1 235,-214 NMOS
M$38 9 21 21 9 NMOS L=1U W=20U AS=40P AD=40P PS=44U PD=44U
* device instance $39 m90 *1 226.5,-214 NMOS
M$39 9 21 7 9 NMOS L=1U W=20U AS=40P AD=40P PS=44U PD=44U
* device instance $40 r180 *1 249,-214 PMOS
M$40 5 5 5 9 PMOS L=1U W=20U AS=40P AD=40P PS=44U PD=44U
* device instance $41 r180 *1 278.5,-143.5 PMOS
M$41 1 10 11 8 PMOS L=1U W=20U AS=40P AD=40P PS=44U PD=44U
* device instance $42 r180 *1 203.5,-144 PMOS
M$42 3 10 18 8 PMOS L=1U W=20U AS=40P AD=40P PS=44U PD=44U
* device instance $43 r180 *1 212.5,-144 PMOS
M$43 3 10 17 8 PMOS L=1U W=20U AS=40P AD=40P PS=44U PD=44U
* device instance $44 r180 *1 225.5,-143.5 PMOS
M$44 6 10 16 8 PMOS L=1U W=20U AS=40P AD=40P PS=44U PD=44U
* device instance $45 r180 *1 234.5,-143.5 PMOS
M$45 6 10 15 8 PMOS L=1U W=20U AS=40P AD=40P PS=44U PD=44U
* device instance $46 r180 *1 247.5,-143.5 PMOS
M$46 5 10 12 8 PMOS L=1U W=20U AS=40P AD=40P PS=44U PD=44U
* device instance $47 r180 *1 256.5,-143.5 PMOS
M$47 5 10 13 8 PMOS L=1U W=20U AS=40P AD=40P PS=44U PD=44U
* device instance $48 r180 *1 269.5,-143.5 PMOS
M$48 1 10 14 8 PMOS L=1U W=20U AS=40P AD=40P PS=44U PD=44U
* device instance $49 m90 *1 236,-185 PMOS
M$49 6 5 21 6 PMOS L=1U W=20U AS=40P AD=40P PS=44U PD=44U
* device instance $50 r0 *1 222.5,-185 PMOS
M$50 6 1 7 6 PMOS L=1U W=20U AS=40P AD=40P PS=44U PD=44U
.ENDS tsd_2021
